LIBRARY ieee;
USE ieee.std_logic_1164.all ;

ENTITY instruction_mem IS
	GENERIC ( N : INTEGER := 32 ) ; 
	PORT ( instruction_mem_address:  IN STD_LOGIC_VECTOR (N-1 DOWNTO 0);
		   instruction: OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0));
END instruction_mem;

ARCHITECTURE Behavior OF instruction_mem IS
BEGIN
	PROCESS (instruction_mem_address)
	BEGIN
		CASE instruction_mem_address IS  -- HERE WE SHOULD HAVE AT LEAST 1 EXAMPLE OF EACH INSTRUCTION IN THE INSTRUCTION SET
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
			WHEN "00000000111111110000000011111111" =>
				instruction <= "00000000111111110000000011111111";
		END CASE;
	END PROCESS;
END Behavior;